module game_control (






);